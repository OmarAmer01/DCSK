/*
================================================================================
* Ring Oscillator With Signal Tap Trigger.
* Author: Omar Tarek Amer
* Date: 12/13/2023
=================================================================================
*/

module ro_sig_tap(
    input i_clk,
    input i_arst_n,
    output o_rand
);

endmodule
