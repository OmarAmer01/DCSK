/*
================================================================================
* Modulator Top Module.
* This module serialls modulates a message with a chaos bit.

* Authors: Omar Tarek Amer

* Date: 12/07/2023
=================================================================================
*/

package spreading_factors_pkg;
  typedef enum {
    SF4  = 0,
    SF8  = 1,
    SF16 = 2,
    SF32 = 3
  } sf_t;
endpackage
