// 3ee4 ya darwee4
//hohoho
