/*
================================================================================
* Modulator Top Module.
* This module serialls modulates a message with a chaos bit.

* Authors: Omar Tarek Amer

* Date: 12/07/2023
=================================================================================
*/

package spreading_factors_pkg;
typedef enum {SF2  = 0,
              SF4  = 1,
              SF8  = 2,
              SF16 = 3} sf_t;
endpackage
